library verilog;
use verilog.vl_types.all;
entity A3_vlg_vec_tst is
end A3_vlg_vec_tst;
