library verilog;
use verilog.vl_types.all;
entity A4_vlg_vec_tst is
end A4_vlg_vec_tst;
