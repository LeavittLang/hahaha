library verilog;
use verilog.vl_types.all;
entity A2ADD16b_vlg_vec_tst is
end A2ADD16b_vlg_vec_tst;
