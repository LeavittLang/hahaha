library verilog;
use verilog.vl_types.all;
entity shift_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        D               : in     vl_logic_vector(15 downto 0);
        GN              : in     vl_logic;
        LR              : in     vl_logic;
        S               : in     vl_logic_vector(1 downto 0);
        sampler_tx      : out    vl_logic
    );
end shift_vlg_sample_tst;
