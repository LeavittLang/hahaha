library verilog;
use verilog.vl_types.all;
entity Atest_vlg_vec_tst is
end Atest_vlg_vec_tst;
