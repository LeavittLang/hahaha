library verilog;
use verilog.vl_types.all;
entity A2_vlg_vec_tst is
end A2_vlg_vec_tst;
