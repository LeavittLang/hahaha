library verilog;
use verilog.vl_types.all;
entity Bus_Latch_vlg_vec_tst is
end Bus_Latch_vlg_vec_tst;
