library verilog;
use verilog.vl_types.all;
entity shift_vlg_vec_tst is
end shift_vlg_vec_tst;
