library verilog;
use verilog.vl_types.all;
entity A_vlg_vec_tst is
end A_vlg_vec_tst;
